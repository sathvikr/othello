module er();

endmodule