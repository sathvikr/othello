module board_manager();

endmodule