module board_manager();

